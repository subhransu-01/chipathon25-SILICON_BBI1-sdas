magic
tech gf180mcuD
timestamp 1755623585
<< nwell >>
rect -18 63 96 127
<< nmos >>
rect 2 21 8 38
rect 19 21 25 38
rect 36 21 42 38
rect 53 21 59 38
rect 70 21 76 38
<< pmos >>
rect 2 72 8 106
rect 19 72 25 106
rect 36 72 42 106
rect 53 72 59 106
rect 70 72 76 106
<< ndiff >>
rect -9 28 2 38
rect -9 23 -6 28
rect -1 23 2 28
rect -9 21 2 23
rect 8 28 19 38
rect 8 23 11 28
rect 16 23 19 28
rect 8 21 19 23
rect 25 28 36 38
rect 25 23 28 28
rect 33 23 36 28
rect 25 21 36 23
rect 42 28 53 38
rect 42 23 45 28
rect 50 23 53 28
rect 42 21 53 23
rect 59 28 70 38
rect 59 23 62 28
rect 67 23 70 28
rect 59 21 70 23
rect 76 28 87 38
rect 76 23 79 28
rect 84 23 87 28
rect 76 21 87 23
<< pdiff >>
rect -9 104 2 106
rect -9 94 -6 104
rect -1 94 2 104
rect -9 72 2 94
rect 8 104 19 106
rect 8 94 11 104
rect 16 94 19 104
rect 8 72 19 94
rect 25 104 36 106
rect 25 94 28 104
rect 33 94 36 104
rect 25 72 36 94
rect 42 104 53 106
rect 42 94 45 104
rect 50 94 53 104
rect 42 72 53 94
rect 59 104 70 106
rect 59 94 62 104
rect 67 94 70 104
rect 59 72 70 94
rect 76 104 87 106
rect 76 94 79 104
rect 84 94 87 104
rect 76 72 87 94
<< ndiffc >>
rect -6 23 -1 28
rect 11 23 16 28
rect 28 23 33 28
rect 45 23 50 28
rect 62 23 67 28
rect 79 23 84 28
<< pdiffc >>
rect -6 94 -1 104
rect 11 94 16 104
rect 28 94 33 104
rect 45 94 50 104
rect 62 94 67 104
rect 79 94 84 104
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 40 12 55 14
rect 40 7 45 12
rect 50 7 55 12
rect 40 5 55 7
rect 74 12 89 14
rect 74 7 79 12
rect 84 7 89 12
rect 74 5 89 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 40 120 56 122
rect 40 115 45 120
rect 50 115 56 120
rect 40 113 56 115
rect 74 120 90 122
rect 74 115 79 120
rect 84 115 90 120
rect 74 113 90 115
<< psubdiffcont >>
rect 11 7 16 12
rect 45 7 50 12
rect 79 7 84 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 45 115 50 120
rect 79 115 84 120
<< polysilicon >>
rect 2 106 8 111
rect 19 106 25 111
rect 36 106 42 111
rect 53 106 59 111
rect 70 106 76 111
rect 2 70 8 72
rect -4 68 8 70
rect -4 62 -2 68
rect 4 62 8 68
rect -4 60 8 62
rect 2 38 8 60
rect 19 70 25 72
rect 19 68 31 70
rect 19 62 23 68
rect 29 62 31 68
rect 19 60 31 62
rect 19 38 25 60
rect 36 51 42 72
rect 53 70 59 72
rect 47 68 59 70
rect 70 68 76 72
rect 47 62 49 68
rect 55 62 76 68
rect 47 60 59 62
rect 30 49 42 51
rect 30 43 32 49
rect 38 43 42 49
rect 30 41 42 43
rect 36 38 42 41
rect 53 38 59 60
rect 70 38 76 62
rect 2 16 8 21
rect 19 16 25 21
rect 36 16 42 21
rect 53 16 59 21
rect 70 16 76 21
<< polycontact >>
rect -2 62 4 68
rect 23 62 29 68
rect 49 62 55 68
rect 32 43 38 49
<< metal1 >>
rect -18 120 96 127
rect -18 115 11 120
rect 16 115 45 120
rect 50 115 79 120
rect 84 115 96 120
rect -18 113 96 115
rect -6 104 -1 106
rect -6 84 -1 94
rect 11 104 16 113
rect 11 92 16 94
rect 28 104 33 106
rect 28 84 33 94
rect 45 104 50 113
rect 45 92 50 94
rect 62 104 67 106
rect -6 79 55 84
rect -4 62 -2 68
rect 4 62 6 68
rect 11 50 16 79
rect 49 68 55 79
rect 21 62 23 68
rect 29 62 31 68
rect 49 60 55 62
rect -6 45 16 50
rect 62 49 67 94
rect 79 104 84 113
rect 79 92 84 94
rect -6 28 -1 45
rect 30 43 32 49
rect 38 43 40 49
rect 62 43 70 49
rect 76 43 79 49
rect -6 21 -1 23
rect 11 28 16 35
rect 11 21 16 23
rect 28 28 33 35
rect 28 21 33 23
rect 45 28 50 30
rect 45 14 50 23
rect 62 28 67 43
rect 62 21 67 23
rect 79 28 84 30
rect 79 14 84 23
rect -18 12 96 14
rect -18 7 11 12
rect 16 7 45 12
rect 50 7 79 12
rect 84 7 96 12
rect -18 0 96 7
<< via1 >>
rect -2 62 4 68
rect 23 62 29 68
rect 32 43 38 49
rect 70 43 76 49
<< metal2 >>
rect -4 68 6 69
rect -4 62 -2 68
rect 4 62 6 68
rect -4 61 6 62
rect 21 68 31 69
rect 21 62 23 68
rect 29 62 31 68
rect 21 61 31 62
rect 30 49 40 50
rect 30 43 32 49
rect 38 43 40 49
rect 30 42 40 43
rect 68 49 78 50
rect 68 43 70 49
rect 76 43 78 49
rect 68 42 78 43
<< labels >>
rlabel nsubdiffcont 13 117 13 117 1 VDD
rlabel psubdiffcont 13 10 13 10 1 VSS
flabel psubdiffcont 11 7 16 12 0 FreeSans 16 0 0 0 VSS
flabel nsubdiffcont 11 115 16 120 0 FreeSans 16 0 0 0 VDD
flabel via1 70 43 76 49 0 FreeSans 32 0 0 0 Y
rlabel nsubdiffcont 45 115 50 120 1 VDD
rlabel nsubdiffcont 79 115 84 120 1 VDD
rlabel psubdiffcont 45 7 50 12 1 VSS
rlabel psubdiffcont 79 7 84 12 1 VSS
flabel pdiffc -6 94 -1 104 0 FreeSans 16 0 0 0 net1
flabel ndiffc 11 23 16 28 0 FreeSans 16 0 0 0 net2
flabel ndiffc 28 23 33 28 0 FreeSans 16 0 0 0 net3
flabel metal2 -2 62 4 68 0 FreeSans 16 0 0 0 A
flabel metal2 23 62 29 68 0 FreeSans 16 0 0 0 B
flabel metal2 32 43 38 49 0 FreeSans 16 0 0 0 C
<< end >>
