magic
tech gf180mcuD
magscale 1 5
timestamp 1755203424
<< error_p >>
rect 52 285 128 293
rect 65 230 75 239
rect 65 220 79 230
<< nwell >>
rect -90 315 535 635
rect 440 310 535 315
<< nmos >>
rect 25 105 55 190
rect 110 105 140 190
rect 165 105 195 190
rect 285 105 315 190
rect 370 105 400 190
<< pmos >>
rect 10 360 40 530
rect 95 360 125 530
rect 180 360 210 530
rect 285 360 315 530
rect 370 360 400 530
<< ndiff >>
rect -45 105 25 190
rect 55 140 110 190
rect 55 115 70 140
rect 95 115 110 140
rect 55 105 110 115
rect 140 105 165 190
rect 195 180 285 190
rect 195 115 210 180
rect 270 115 285 180
rect 195 105 285 115
rect 315 140 370 190
rect 315 115 330 140
rect 355 115 370 140
rect 315 105 370 115
rect 400 140 455 190
rect 400 115 415 140
rect 440 115 455 140
rect 400 105 455 115
<< pdiff >>
rect -45 520 10 530
rect -45 370 -30 520
rect -5 370 10 520
rect -45 360 10 370
rect 40 520 95 530
rect 40 370 55 520
rect 80 370 95 520
rect 40 360 95 370
rect 125 520 180 530
rect 125 370 140 520
rect 165 370 180 520
rect 125 360 180 370
rect 210 520 285 530
rect 210 370 225 520
rect 270 370 285 520
rect 210 360 285 370
rect 315 520 370 530
rect 315 470 330 520
rect 355 470 370 520
rect 315 360 370 470
rect 400 520 455 530
rect 400 470 415 520
rect 440 470 455 520
rect 400 360 455 470
<< ndiffc >>
rect 70 115 95 140
rect 210 115 270 180
rect 330 115 355 140
rect 415 115 440 140
<< pdiffc >>
rect -30 370 -5 520
rect 55 370 80 520
rect 140 370 165 520
rect 225 370 270 520
rect 330 470 355 520
rect 415 470 440 520
<< psubdiff >>
rect 30 60 105 70
rect 30 35 55 60
rect 80 35 105 60
rect 30 25 105 35
rect 150 60 225 70
rect 150 35 175 60
rect 200 35 225 60
rect 150 25 225 35
rect 270 60 345 70
rect 270 35 295 60
rect 320 35 345 60
rect 270 25 345 35
<< nsubdiff >>
rect 30 600 105 610
rect 30 575 55 600
rect 80 575 105 600
rect 30 565 105 575
rect 150 600 225 610
rect 150 575 175 600
rect 200 575 225 600
rect 150 565 225 575
rect 270 600 345 610
rect 270 575 295 600
rect 320 575 345 600
rect 270 565 345 575
<< psubdiffcont >>
rect 55 35 80 60
rect 175 35 200 60
rect 295 35 320 60
<< nsubdiffcont >>
rect 55 575 80 600
rect 175 575 200 600
rect 295 575 320 600
<< polysilicon >>
rect 10 530 40 555
rect 95 530 125 555
rect 180 530 210 555
rect 285 530 315 555
rect 370 530 400 555
rect 10 255 40 360
rect 95 270 125 360
rect 180 335 210 360
rect 180 325 245 335
rect 180 315 205 325
rect -30 245 40 255
rect -30 215 -20 245
rect 10 215 40 245
rect 65 260 125 270
rect 65 230 75 260
rect 105 230 125 260
rect 165 295 205 315
rect 235 295 245 325
rect 165 285 245 295
rect 65 220 140 230
rect -30 205 55 215
rect 25 190 55 205
rect 110 190 140 220
rect 165 190 195 285
rect 285 270 315 360
rect 265 260 315 270
rect 265 230 275 260
rect 305 230 315 260
rect 265 220 315 230
rect 285 190 315 220
rect 370 190 400 360
rect 25 80 55 105
rect 110 80 140 105
rect 165 80 195 105
rect 285 80 315 105
rect 370 80 400 105
<< polycontact >>
rect -20 215 10 245
rect 75 230 105 260
rect 205 295 235 325
rect 275 230 305 260
<< metal1 >>
rect -90 600 535 635
rect -90 575 55 600
rect 80 575 175 600
rect 200 575 295 600
rect 320 575 535 600
rect -90 565 535 575
rect -30 520 -5 530
rect -30 310 -5 370
rect 55 520 80 565
rect 55 360 80 370
rect 140 520 165 530
rect 140 310 165 370
rect 225 520 270 565
rect 225 360 270 370
rect 330 520 355 530
rect 330 335 355 470
rect 415 520 440 530
rect 415 335 440 470
rect -30 285 165 310
rect 195 295 205 325
rect 235 295 245 325
rect 330 310 440 335
rect 75 260 105 270
rect -20 245 10 255
rect 75 220 105 230
rect 140 260 165 285
rect 275 260 305 270
rect 140 230 275 260
rect -20 205 10 215
rect 140 180 165 230
rect 275 220 305 230
rect 70 155 165 180
rect 210 180 270 190
rect 70 140 95 155
rect 70 105 95 115
rect 210 70 270 115
rect 330 140 355 310
rect 330 105 355 115
rect 415 280 440 310
rect 415 250 450 280
rect 480 250 490 280
rect 415 140 440 250
rect 415 105 440 115
rect -90 60 535 70
rect -90 35 55 60
rect 80 35 175 60
rect 200 35 295 60
rect 320 35 535 60
rect -90 0 535 35
<< via1 >>
rect 205 295 235 325
rect -20 215 10 245
rect 75 230 105 260
rect 450 250 480 280
<< metal2 >>
rect 195 325 245 330
rect 195 295 205 325
rect 235 295 245 325
rect 195 290 245 295
rect 445 280 485 285
rect 65 260 120 270
rect -30 245 20 255
rect -30 215 -20 245
rect 10 215 20 245
rect 65 230 75 260
rect 105 230 120 260
rect 445 250 450 280
rect 480 250 485 280
rect 445 245 485 250
rect 65 220 120 230
rect -30 205 20 215
<< labels >>
rlabel nsubdiffcont 65 585 65 585 1 VDD
rlabel psubdiffcont 65 50 65 50 1 VSS
flabel psubdiffcont 55 35 80 60 0 FreeSans 80 0 0 0 VSS
flabel nsubdiffcont 55 575 80 600 0 FreeSans 80 0 0 0 VDD
flabel via1 450 250 480 280 0 FreeSans 160 0 0 0 Y
flabel metal2 205 295 235 325 0 FreeSans 160 0 0 0 C
flabel metal2 -20 215 10 245 0 FreeSans 160 0 0 0 A
flabel metal2 75 230 105 260 0 FreeSans 160 0 0 0 B
<< end >>
