magic
tech gf180mcuD
timestamp 1755257249
<< nwell >>
rect -18 63 94 127
<< nmos >>
rect 5 21 11 38
rect 22 21 28 38
rect 33 21 39 38
rect 57 21 63 38
rect 74 21 80 38
<< pmos >>
rect 2 72 8 106
rect 19 72 25 106
rect 36 72 42 106
rect 57 72 63 106
rect 74 72 80 106
<< ndiff >>
rect -9 28 5 38
rect -9 23 -3 28
rect 2 23 5 28
rect -9 21 5 23
rect 11 21 22 38
rect 28 21 33 38
rect 39 36 57 38
rect 39 23 42 36
rect 54 23 57 36
rect 39 21 57 23
rect 63 28 74 38
rect 63 23 66 28
rect 71 23 74 28
rect 63 21 74 23
rect 80 21 85 38
<< pdiff >>
rect -9 104 2 106
rect -9 74 -6 104
rect -1 74 2 104
rect -9 72 2 74
rect 8 104 19 106
rect 8 74 11 104
rect 16 74 19 104
rect 8 72 19 74
rect 25 104 36 106
rect 25 74 28 104
rect 33 74 36 104
rect 25 72 36 74
rect 42 104 57 106
rect 42 74 45 104
rect 54 74 57 104
rect 42 72 57 74
rect 63 104 74 106
rect 63 94 66 104
rect 71 94 74 104
rect 63 72 74 94
rect 80 72 85 106
<< ndiffc >>
rect -3 23 2 28
rect 42 23 54 36
rect 66 23 71 28
<< pdiffc >>
rect -6 74 -1 104
rect 11 74 16 104
rect 28 74 33 104
rect 45 74 54 104
rect 66 94 71 104
<< psubdiff >>
rect 6 12 21 14
rect 6 7 11 12
rect 16 7 21 12
rect 6 5 21 7
rect 30 12 45 14
rect 30 7 35 12
rect 40 7 45 12
rect 30 5 45 7
rect 54 12 69 14
rect 54 7 59 12
rect 64 7 69 12
rect 54 5 69 7
<< nsubdiff >>
rect 6 120 21 122
rect 6 115 11 120
rect 16 115 21 120
rect 6 113 21 115
rect 30 120 45 122
rect 30 115 35 120
rect 40 115 45 120
rect 30 113 45 115
rect 54 120 69 122
rect 54 115 59 120
rect 64 115 69 120
rect 54 113 69 115
<< psubdiffcont >>
rect 11 7 16 12
rect 35 7 40 12
rect 59 7 64 12
<< nsubdiffcont >>
rect 11 115 16 120
rect 35 115 40 120
rect 59 115 64 120
<< polysilicon >>
rect 2 106 8 111
rect 19 106 25 111
rect 36 106 42 111
rect 57 106 63 111
rect 74 106 80 111
rect 2 53 8 72
rect 19 58 25 72
rect 36 67 42 72
rect 57 69 63 72
rect 74 69 80 72
rect 36 65 49 67
rect 36 63 41 65
rect -8 50 8 53
rect -8 44 -5 50
rect 1 44 8 50
rect 13 56 25 58
rect 13 50 15 56
rect 21 52 25 56
rect 33 59 41 63
rect 47 59 49 65
rect 33 57 49 59
rect 57 63 80 69
rect 21 50 26 52
rect 13 49 26 50
rect 14 48 26 49
rect 22 47 26 48
rect -8 41 11 44
rect 5 38 11 41
rect 22 38 28 47
rect 33 38 39 57
rect 57 54 63 63
rect 53 52 63 54
rect 53 46 55 52
rect 61 47 63 52
rect 74 47 80 63
rect 61 46 80 47
rect 53 44 80 46
rect 57 41 80 44
rect 57 38 63 41
rect 74 38 80 41
rect 5 16 11 21
rect 22 16 28 21
rect 33 16 39 21
rect 57 16 63 21
rect 74 16 80 21
<< polycontact >>
rect -5 44 1 50
rect 15 50 21 56
rect 41 59 47 65
rect 55 46 61 52
<< metal1 >>
rect -18 120 94 127
rect -18 115 11 120
rect 16 115 35 120
rect 40 115 59 120
rect 64 115 94 120
rect -18 113 94 115
rect -6 104 -1 106
rect -6 67 -1 74
rect 11 104 16 113
rect 11 72 16 74
rect 28 104 33 106
rect 28 67 33 74
rect 45 104 54 113
rect 45 72 54 74
rect 66 104 71 106
rect -6 62 33 67
rect 13 50 15 56
rect 21 50 23 56
rect 28 52 33 62
rect 39 59 41 65
rect 47 59 49 65
rect 66 59 71 94
rect 55 52 61 54
rect -7 44 -5 50
rect 1 44 3 50
rect 28 46 55 52
rect 28 36 33 46
rect 55 44 61 46
rect 66 53 73 59
rect 79 53 81 59
rect -3 31 33 36
rect 42 36 54 38
rect -3 28 2 31
rect -3 21 2 23
rect 42 14 54 23
rect 66 28 71 53
rect 66 21 71 23
rect -18 12 94 14
rect -18 7 11 12
rect 16 7 35 12
rect 40 7 59 12
rect 64 7 94 12
rect -18 0 94 7
<< via1 >>
rect 15 50 21 56
rect 41 59 47 65
rect -5 44 1 50
rect 73 53 79 59
<< metal2 >>
rect 39 65 49 66
rect 39 59 41 65
rect 47 59 49 65
rect 39 58 49 59
rect 72 59 80 60
rect 13 56 23 57
rect -7 50 3 51
rect -7 44 -5 50
rect 1 44 3 50
rect 13 50 15 56
rect 21 50 23 56
rect 72 53 73 59
rect 79 53 80 59
rect 72 52 80 53
rect 13 49 23 50
rect -7 43 3 44
<< labels >>
rlabel nsubdiffcont 13 117 13 117 1 VDD
rlabel psubdiffcont 13 10 13 10 1 VSS
flabel psubdiffcont 11 7 16 12 0 FreeSans 16 0 0 0 VSS
flabel nsubdiffcont 11 115 16 120 0 FreeSans 16 0 0 0 VDD
flabel metal2 41 59 47 65 0 FreeSans 32 0 0 0 C
flabel metal2 -5 44 1 50 0 FreeSans 32 0 0 0 A
flabel metal2 15 50 21 56 0 FreeSans 32 0 0 0 B
flabel via1 73 53 79 59 0 FreeSans 32 0 0 0 Y
<< end >>
