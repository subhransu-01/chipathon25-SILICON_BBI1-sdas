magic
tech gf180mcuD
timestamp 1756608592
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_0
timestamp 1756569562
transform 1 0 17 0 1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_1
timestamp 1756569562
transform 1 0 17 0 -1 332
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_2
timestamp 1756569562
transform 1 0 17 0 -1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_3
timestamp 1756569562
transform 1 0 95 0 -1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_4
timestamp 1756569562
transform 1 0 173 0 -1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_5
timestamp 1756569562
transform 1 0 251 0 -1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_6
timestamp 1756569562
transform 1 0 95 0 1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_7
timestamp 1756569562
transform 1 0 173 0 1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_8
timestamp 1756569562
transform 1 0 251 0 1 0
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_9
timestamp 1756569562
transform 1 0 95 0 -1 332
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_10
timestamp 1756569562
transform 1 0 173 0 -1 332
box -17 0 61 166
use gf180mcu_osu_sc_gp12t3v3__nand3_1  gf180mcu_osu_sc_gp12t3v3__nand3_1_11
timestamp 1756569562
transform 1 0 251 0 -1 332
box -17 0 61 166
<< end >>
