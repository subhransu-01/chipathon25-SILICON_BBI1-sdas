magic
tech gf180mcuD
timestamp 1756607006
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_0
timestamp 1756568175
transform 1 0 -114 0 1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_1
timestamp 1756568175
transform 1 0 -36 0 1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_2
timestamp 1756568175
transform 1 0 42 0 1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_3
timestamp 1756568175
transform 1 0 -192 0 1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_4
timestamp 1756568175
transform 1 0 -192 0 -1 254
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_5
timestamp 1756568175
transform 1 0 -114 0 -1 254
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_6
timestamp 1756568175
transform 1 0 -36 0 -1 254
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_7
timestamp 1756568175
transform 1 0 42 0 -1 254
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_8
timestamp 1756568175
transform 1 0 -192 0 -1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_9
timestamp 1756568175
transform 1 0 -114 0 -1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_10
timestamp 1756568175
transform 1 0 -36 0 -1 0
box 114 0 192 127
use gf180mcu_osu_sc_gp9t3v3__nor3_1  gf180mcu_osu_sc_gp9t3v3__nor3_1_11
timestamp 1756568175
transform 1 0 42 0 -1 0
box 114 0 192 127
<< end >>
