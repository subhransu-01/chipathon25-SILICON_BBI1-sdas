magic
tech gf180mcuD
timestamp 1755641212
<< nwell >>
rect 105 63 200 127
<< nmos >>
rect 124 21 130 38
rect 141 21 147 38
rect 158 21 164 38
rect 175 21 181 38
<< pmos >>
rect 124 72 130 106
rect 141 72 147 106
rect 158 72 164 106
rect 175 72 181 106
<< ndiff >>
rect 114 29 124 38
rect 114 23 116 29
rect 121 23 124 29
rect 114 21 124 23
rect 130 29 141 38
rect 130 23 133 29
rect 138 23 141 29
rect 130 21 141 23
rect 147 29 158 38
rect 147 23 150 29
rect 155 23 158 29
rect 147 21 158 23
rect 164 29 175 38
rect 164 23 167 29
rect 172 23 175 29
rect 164 21 175 23
rect 181 29 191 38
rect 181 23 184 29
rect 189 23 191 29
rect 181 21 191 23
<< pdiff >>
rect 114 104 124 106
rect 114 90 116 104
rect 121 90 124 104
rect 114 72 124 90
rect 130 104 141 106
rect 130 90 133 104
rect 138 90 141 104
rect 130 72 141 90
rect 147 104 158 106
rect 147 90 150 104
rect 155 90 158 104
rect 147 72 158 90
rect 164 104 175 106
rect 164 90 167 104
rect 172 90 175 104
rect 164 72 175 90
rect 181 104 191 106
rect 181 90 184 104
rect 189 90 191 104
rect 181 72 191 90
<< ndiffc >>
rect 116 23 121 29
rect 133 23 138 29
rect 150 23 155 29
rect 167 23 172 29
rect 184 23 189 29
<< pdiffc >>
rect 116 90 121 104
rect 133 90 138 104
rect 150 90 155 104
rect 167 90 172 104
rect 184 90 189 104
<< psubdiff >>
rect 111 12 126 14
rect 111 7 116 12
rect 121 7 126 12
rect 111 5 126 7
rect 145 12 160 14
rect 145 7 150 12
rect 155 7 160 12
rect 145 5 160 7
rect 179 12 194 14
rect 179 7 184 12
rect 189 7 194 12
rect 179 5 194 7
<< nsubdiff >>
rect 111 120 126 122
rect 111 115 116 120
rect 121 115 126 120
rect 111 113 126 115
rect 145 120 160 122
rect 145 115 150 120
rect 155 115 160 120
rect 145 113 160 115
rect 179 120 194 122
rect 179 115 185 120
rect 190 115 194 120
rect 179 113 194 115
<< psubdiffcont >>
rect 116 7 121 12
rect 150 7 155 12
rect 184 7 189 12
<< nsubdiffcont >>
rect 116 115 121 120
rect 150 115 155 120
rect 185 115 190 120
<< polysilicon >>
rect 124 106 130 111
rect 141 106 147 111
rect 158 106 164 111
rect 175 106 181 111
rect 124 70 130 72
rect 118 68 130 70
rect 118 62 120 68
rect 126 62 130 68
rect 118 60 130 62
rect 124 38 130 60
rect 141 70 147 72
rect 141 68 153 70
rect 141 62 145 68
rect 151 62 153 68
rect 141 60 153 62
rect 141 38 147 60
rect 158 50 164 72
rect 175 70 181 72
rect 169 68 181 70
rect 169 62 171 68
rect 177 62 181 68
rect 169 60 181 62
rect 158 48 170 50
rect 158 42 162 48
rect 168 42 170 48
rect 158 40 170 42
rect 158 38 164 40
rect 175 38 181 60
rect 124 16 130 21
rect 141 16 147 21
rect 158 16 164 21
rect 175 16 181 21
<< polycontact >>
rect 120 62 126 68
rect 145 62 151 68
rect 171 62 177 68
rect 162 42 168 48
<< metal1 >>
rect 105 120 200 127
rect 105 115 116 120
rect 121 115 150 120
rect 155 115 185 120
rect 190 115 200 120
rect 105 113 200 115
rect 116 104 121 106
rect 116 81 121 90
rect 133 104 138 106
rect 133 88 138 90
rect 150 104 155 106
rect 150 88 155 90
rect 167 104 172 113
rect 167 88 172 90
rect 184 104 189 106
rect 116 76 177 81
rect 118 62 120 68
rect 126 62 128 68
rect 133 41 138 76
rect 171 68 177 76
rect 143 62 145 68
rect 151 62 153 68
rect 171 60 177 62
rect 160 42 162 48
rect 168 42 170 48
rect 184 47 189 90
rect 184 41 190 47
rect 196 41 198 47
rect 116 36 155 41
rect 116 29 121 36
rect 116 21 121 23
rect 133 29 138 31
rect 133 14 138 23
rect 150 29 155 36
rect 150 21 155 23
rect 167 29 172 31
rect 150 14 155 15
rect 167 14 172 23
rect 184 29 189 41
rect 184 21 189 23
rect 105 12 200 14
rect 105 7 116 12
rect 121 7 150 12
rect 155 7 184 12
rect 189 7 200 12
rect 105 0 200 7
<< via1 >>
rect 120 62 126 68
rect 145 62 151 68
rect 162 42 168 48
rect 190 41 196 47
<< metal2 >>
rect 118 68 128 69
rect 118 62 120 68
rect 126 62 128 68
rect 118 61 128 62
rect 143 68 153 69
rect 143 62 145 68
rect 151 62 153 68
rect 143 61 153 62
rect 160 48 170 49
rect 160 42 162 48
rect 168 42 170 48
rect 160 41 170 42
rect 188 47 198 48
rect 188 41 190 47
rect 196 41 198 47
rect 188 40 198 41
<< labels >>
rlabel nsubdiffcont 116 115 121 120 1 VDD
rlabel nsubdiffcont 150 115 155 120 1 VDD
rlabel nsubdiffcont 185 115 190 120 1 VDD
rlabel psubdiffcont 116 7 121 12 1 VSS
rlabel psubdiffcont 150 7 155 12 1 VSS
rlabel psubdiffcont 184 7 189 12 1 VSS
rlabel metal2 120 62 126 68 1 A
rlabel metal2 145 62 151 68 1 B
rlabel via1 190 41 196 47 1 Y
rlabel metal2 162 42 168 48 1 C
rlabel pdiffc 133 90 138 104 1 net2
rlabel ndiffc 116 23 121 29 1 net3
rlabel pdiffc 150 90 155 104 1 net1
<< end >>
