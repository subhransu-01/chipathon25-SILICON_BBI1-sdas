magic
tech gf180mcuD
magscale 1 10
timestamp 1755148472
<< error_p >>
rect -99 140 -90 169
rect -70 60 -61 140
rect 0 60 9 169
rect 160 50 169 169
rect 350 -250 400 -244
rect 350 -263 393 -250
rect 350 -277 363 -263
rect 350 -290 393 -277
rect -200 -373 -140 -354
rect -200 -387 -187 -373
rect 50 -383 120 -370
rect 210 -383 260 -370
rect -200 -400 -140 -387
rect -296 -410 -130 -404
rect 107 -407 120 -383
rect 247 -407 260 -383
rect 50 -420 120 -407
rect 210 -420 260 -407
<< nwell >>
rect -430 460 590 470
rect -430 -190 760 460
<< nmos >>
rect -150 -650 -90 -520
rect 0 -650 60 -520
rect 160 -650 220 -520
rect 380 -650 440 -520
<< pmos >>
rect -150 30 -90 160
rect 0 30 60 160
rect 160 30 220 160
rect 380 30 440 160
<< ndiff >>
rect -260 -540 -150 -520
rect -260 -610 -240 -540
rect -190 -610 -150 -540
rect -260 -650 -150 -610
rect -90 -650 0 -520
rect 60 -650 160 -520
rect 220 -560 380 -520
rect 220 -630 250 -560
rect 350 -630 380 -560
rect 220 -650 380 -630
rect 440 -650 630 -520
<< pdiff >>
rect -110 320 20 340
rect -110 250 -90 320
rect 0 250 20 320
rect -110 230 20 250
rect 230 320 370 340
rect 230 250 250 320
rect 350 250 370 320
rect 230 230 370 250
rect -260 140 -150 160
rect -260 50 -240 140
rect -190 50 -150 140
rect -260 30 -150 50
rect -90 140 0 160
rect -90 60 -70 140
rect -20 60 0 140
rect -90 30 0 60
rect 60 140 160 160
rect 60 50 90 140
rect 140 50 160 140
rect 60 30 160 50
rect 220 140 380 160
rect 220 60 250 140
rect 350 60 380 140
rect 220 30 380 60
rect 440 30 630 160
rect 210 -820 390 -800
rect 210 -870 240 -820
rect 360 -870 390 -820
rect 210 -890 390 -870
<< ndiffc >>
rect -240 -610 -190 -540
rect 250 -630 350 -560
<< pdiffc >>
rect -90 250 0 320
rect 250 250 350 320
rect -240 50 -190 140
rect -70 60 -20 140
rect 90 50 140 140
rect 250 60 350 140
rect 240 -870 360 -820
<< polysilicon >>
rect -150 160 -90 210
rect 0 160 60 210
rect 160 160 220 210
rect 380 160 440 210
rect -150 -360 -90 30
rect -140 -400 -90 -360
rect -150 -520 -90 -400
rect 0 -370 60 30
rect 160 -370 220 30
rect 380 -250 440 30
rect 400 -290 440 -250
rect 0 -420 50 -370
rect 160 -420 210 -370
rect 0 -520 60 -420
rect 160 -520 220 -420
rect 380 -520 440 -290
rect -150 -710 -90 -650
rect 0 -710 60 -650
rect 160 -710 220 -650
rect 380 -710 440 -650
<< polycontact >>
rect -200 -400 -140 -360
rect 350 -290 400 -250
rect 50 -420 120 -370
rect 210 -420 260 -370
<< metal1 >>
rect -260 320 500 400
rect -260 250 -90 320
rect 0 250 250 320
rect 350 250 500 320
rect -260 230 500 250
rect -250 140 -150 160
rect -250 50 -240 140
rect -190 50 -150 140
rect -250 30 -150 50
rect -70 140 -20 230
rect -70 40 -20 60
rect 60 140 160 160
rect 60 50 90 140
rect 140 50 160 140
rect 60 30 160 50
rect 240 140 360 230
rect 240 60 250 140
rect 350 60 360 140
rect 240 40 360 60
rect -250 -240 -170 30
rect 70 -240 150 30
rect -250 -250 420 -240
rect -250 -290 350 -250
rect 400 -290 420 -250
rect -250 -300 420 -290
rect 470 -270 610 140
rect -320 -360 -130 -350
rect -320 -400 -200 -360
rect -140 -400 -130 -360
rect -320 -410 -130 -400
rect -80 -450 -10 -300
rect 40 -370 130 -360
rect 40 -420 50 -370
rect 120 -420 130 -370
rect 40 -430 130 -420
rect 190 -370 280 -360
rect 190 -420 210 -370
rect 260 -420 280 -370
rect 190 -430 280 -420
rect 470 -410 670 -270
rect -250 -510 -10 -450
rect -250 -540 -160 -510
rect -250 -610 -240 -540
rect -190 -610 -160 -540
rect -250 -630 -160 -610
rect 230 -560 370 -540
rect 230 -630 250 -560
rect 350 -630 370 -560
rect 470 -630 610 -410
rect 230 -790 370 -630
rect -260 -820 490 -790
rect -260 -870 240 -820
rect 360 -870 490 -820
rect -260 -950 490 -870
<< labels >>
flabel metal1 -80 370 280 370 0 FreeSans 480 0 0 0 VDD
flabel metal1 -160 -930 370 -930 1 FreeSans 480 0 0 0 GND
flabel metal1 -140 -400 -140 -360 7 FreeSans 480 0 0 0 A
flabel metal1 50 -420 50 -370 3 FreeSans 480 0 0 0 B
flabel metal1 210 -420 210 -370 3 FreeSans 480 0 0 0 C
flabel metal1 660 -410 670 -280 7 FreeSans 480 0 0 0 Y
<< end >>
